LIBRARY IEEE;
LIBRARY ALTERA_MF;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ALTERA_MF.ALTERA_MF_COMPONENTS.ALL;
USE LPM.LPM_COMPONENTS.ALL;

--initializes the input/outputs of the state machine
ENTITY SRAM IS
	PORT(
		IO_WRITE    	: IN    STD_LOGIC;
		SRAM_ADHI_EN   	: IN    STD_LOGIC;
		SRAM_ADLOW_EN   : IN    STD_LOGIC;
		SRAM_WRITE	    : IN    STD_LOGIC;
		SRAM_READ   	: IN    STD_LOGIC;
		CLOCK			: IN    STD_LOGIC;          
		IO_DATA  		: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR  		: OUT   STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_OE_N 		: OUT   STD_LOGIC;
		SRAM_DQ			: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_WE_N		: OUT   STD_LOGIC;
		SRAM_UB_N		: OUT   STD_LOGIC;
		SRAM_LB_N		: OUT   STD_LOGIC;
		SRAM_CE_N		: OUT   STD_LOGIC
	);
END SRAM;

ARCHITECTURE a OF SRAM IS

--defines the states of the I/O device
TYPE STATE_TYPE IS (
		IDLE,
		WRITE_EN, 
		DATA_SEND, 
		WRITE_DISABLE,
		READ_DATA1, 
		READ_DATA2, 
		READ_DATA3
	);
--made a signal called state we can can referece this instead of STATE_TYPE
SIGNAL STATE: STATE_TYPE;

BEGIN

--these three all go to ground, so here they are zero
SRAM_UB_N <= '0';
SRAM_LB_N <= '0';
SRAM_CE_N <= '0';

	PROCESS (IO_WRITE, SRAM_ADHI_EN)
	BEGIN
		IF (IO_WRITE = '1') AND (SRAM_ADHI_EN = '1') THEN
			SRAM_ADDR(17 DOWNTO 16) <= IO_DATA(1 DOWNTO 0);
		END IF;
	END PROCESS;

	PROCESS (IO_WRITE, SRAM_ADLOW_EN)	
	BEGIN	
		IF (IO_WRITE = '1') AND (SRAM_ADLOW_EN = '1') THEN
			SRAM_ADDR(15 DOWNTO 0) <= IO_DATA;
		END IF;
	END PROCESS;

	PROCESS (IO_WRITE, CLOCK, SRAM_WRITE, SRAM_READ)
	BEGIN
		IF (IO_WRITE = '0') THEN          
			STATE <= IDLE;
		ELSE IF (RISING_EDGE(CLOCK)) THEN
			CASE STATE IS
				--Write
				WHEN WRITE_EN => 
					SRAM_WE_N <= '0';
					STATE <= DATA_SEND;
				WHEN DATA_SEND =>
					SRAM_DQ <= IO_DATA;
					STATE <= WRITE_DISABLE;
				WHEN WRITE_DISABLE =>
					SRAM_WE_N <= '1';
					IO_DATA <= "ZZZZZZZZZZZZZZZZ";
				--Read
				WHEN READ_DATA1 =>
					SRAM_OE_N <= '0';
					STATE <= READ_DATA2;
				WHEN READ_DATA2 =>
					STATE <= READ_DATA3;
				WHEN READ_DATA3 =>
					IO_DATA <= SRAM_DQ;
					SRAM_OE_N <= '1';
				
	
	END PROCESS;
	
--		
--	
--PROCESS (CLOCK, IO_WRITE, SRAM_WRITE)
--BEGIN 
--	IF (IO_WRITE = '1') AND (SRAM_WRITE = '1') THEN
--		IF (RISING_EDGE(CLOCK)) THEN
--			STATE <= WRITE_EN;
--			CASE STATE IS
--				WHEN WRITE_EN =>
--					SRAM_WE_N <= '0';
--					STATE <= DATA_SEND;
--				WHEN DATA_SEND =>
--					SRAM_DQ <= IO_DATA;
--					STATE <= WRITE_DISABLE;
--				WHEN WRITE_DISABLE =>
--					SRAM_WE_N <= '1';
--					IO_DATA <= "ZZZZZZZZZZZZZZZZ";
--				WHEN OTHERS =>
--			END CASE;
--		END IF;
--	END IF;
--END PROCESS;
--
--
--PROCESS (CLOCK, SRAM_READ, IO_WRITE)
--BEGIN
--	IF (IO_WRITE = '1') AND (SRAM_READ = '1') THEN
--		IF (RISING_EDGE(CLOCK)) THEN
--			STATE <= READ_DATA1;
--			CASE STATE IS
--				WHEN DATA_SEND =>
--					SRAM_DQ <= IO_DATA;
--					STATE <= WRITE_DISABLE;
--				WHEN WRITE_DISABLE =>
--					SRAM_WE_N <= '1';
--					IO_DATA <= "ZZZZZZZZZZZZZZZZ";
--				WHEN OTHERS =>
--			END CASE;
--		END IF;
--	END IF;
--END PROCESS;


























END a;