LIBRARY IEEE;
LIBRARY ALTERA_MF;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ALTERA_MF.ALTERA_MF_COMPONENTS.ALL;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY SRAM IS
	PORT(
		IO_WRITE    	: IN    STD_LOGIC;
		SRAM_ADHI_EN   	: IN    STD_LOGIC;
		SRAM_ADLOW_EN   : IN    STD_LOGIC;
		SRAM_WRITE	    : IN    STD_LOGIC;
		SRAM_READ   	: IN    STD_LOGIC;
		IO_DATA  		: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR  		: OUT   STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_OE_N 		: OUT   STD_LOGIC;
		SRAM_DQ			: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_WE_N		: OUT   STD_LOGIC;
		SRAM_UB_N		: OUT   STD_LOGIC;
		SRAM_LB_N		: OUT   STD_LOGIC;
		SRAM_CE_N		: OUT   STD_LOGIC
	);
END SRAM;

ARCHITECTURE a OF SRAM IS
BEGIN
END a;