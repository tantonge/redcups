LIBRARY IEEE;
LIBRARY ALTERA_MF;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ALTERA_MF.ALTERA_MF_COMPONENTS.ALL;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY SRAM IS
	PORT(
		IO_WRITE    	: IN    STD_LOGIC;
		SRAM_ADHI_EN   	: IN    STD_LOGIC;
		SRAM_ADLOW_EN   : IN    STD_LOGIC;
		SRAM_WRITE	    : IN    STD_LOGIC;
		SRAM_READ   	: IN    STD_LOGIC;
		IO_DATA  		: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR  		: OUT   STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_OE_N 		: OUT   STD_LOGIC;
		SRAM_DQ			: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_WE_N		: OUT   STD_LOGIC;
		SRAM_UB_N		: OUT   STD_LOGIC;
		SRAM_LB_N		: OUT   STD_LOGIC;
		SRAM_CE_N		: OUT   STD_LOGIC
	);
END SRAM;

ARCHITECTURE a OF SRAM IS

TYPE STATE_TYPE IS (
		RESET_PC, FETCH, DECODE
	);
	
BEGIN

SRAM_UB_N <= '0';
SRAM_LB_N <= '0';
SRAM_CE_N <= '0';

PROCESS IS
BEGIN 
SRAM_OE_N <= '1';
SRAM_WE_N <= '1';
WAIT UNTIL (IO_WRITE = '1');
	IF (SRAM_ADHI_EN = '1') THEN
		SRAM_ADDR(17 DOWNTO 16) <= IO_DATA(1 DOWNTO 0);
	END IF;
		
	IF (SRAM_ADLOW_EN = '1') THEN
		SRAM_ADDR(15 DOWNTO 0) <= IO_DATA;
	END IF;
		
	IF (SRAM_WRITE = '1') THEN
		SRAM_WE_N <= '0';
		WAIT FOR 25 ns;
		SRAM_DQ <= IO_DATA;
		WAIT FOR 25 ns;
		SRAM_WE_N <= '1';
		WAIT FOR 1 ns;
		IO_DATA <= "ZZZZZZZZZZZZZZZZ";
	END IF;
	
	IF (SRAM_READ = '1') THEN
		SRAM_OE_N <= '0';
		WAIT FOR 50 ns;
		IO_DATA <= SRAM_DQ;
		WAIT FOR 400 ns;
		SRAM_OE_N <= '1';
	END IF;
	
END PROCESS;

END a;